interface adder();

	logic a_in, b_in, c_in;
	logic carry_out, sum_out;

endinterface
