program helloworld();
	initial begin
		$display("hello world!");
	end



endprogram
