program test();
	initial begin
		$display("tt");
	end



endprogram
